library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RED is
    Port (
        RED_INPUT : in  STD_LOGIC_VECTOR(7 downto 0);
		  RED_CLOCK   : in  STD_LOGIC
	 );
end RED;

architecture Behavioral of RED is
begin


    process(RED_INPUT,RED_CLOCK)
    begin

	 
	 
	 
        null;
    end process;
end Behavioral;
